** Profile: "SCHEMATIC1-JEDL_Project_1"  [ C:\Users\EvanB\Desktop\JEDL_Project_1-master\jedl_project_1-pspicefiles\schematic1\jedl_project_1.sim ] 

** Creating circuit file "JEDL_Project_1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../jedl_project_1-pspicefiles/jedl_project_1.lib" 
* From [PSPICE NETLIST] section of C:\SPB_DATA\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 0.6 0 0.001 SKIPBP 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
